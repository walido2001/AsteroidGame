module main(input hello, output bye);

endmodule